VHDL