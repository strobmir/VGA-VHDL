VHDL

VHDL2